// tb_myproject_inst.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module tb_myproject_inst (
		input  wire          start,      //       call.valid
		output wire          busy,       //           .stall
		input  wire          clock,      //      clock.clk
		input  wire [3135:0] inputs,     //     inputs.data
		input  wire          resetn,     //      reset.reset_n
		output wire          done,       //     return.valid
		input  wire          stall,      //           .stall
		output wire [159:0]  returndata  // returndata.data
	);

	myproject_internal myproject_internal_inst (
		.clock      (clock),      //      clock.clk
		.resetn     (resetn),     //      reset.reset_n
		.start      (start),      //       call.valid
		.busy       (busy),       //           .stall
		.done       (done),       //     return.valid
		.stall      (stall),      //           .stall
		.returndata (returndata), // returndata.data
		.inputs     (inputs)      //     inputs.data
	);

endmodule
